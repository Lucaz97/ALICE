`timescale 1ns / 1ps

module c_mod(a, b, c);

input a, c;
output b; 

assign b = a; 

endmodule 