

module b_mod(in1, out1);



input in1;
output out1; 


c_mod	c_inst0(
		.a(	in1	),
		.b(	out1 )
		);

 
endmodule 