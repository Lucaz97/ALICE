
module a_mod(in1, out1);


input in1;
output out1; 


b_mod	b_inst0(
		.in1(	in1	),
		.out1(	out1		)
		);

endmodule